LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		endereco : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saida : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE arranjo_memoria IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(19 DOWNTO 0);
	
	-- para ganhar: R L D R
															--	R	U	L	D
	SIGNAL memoria : arranjo_memoria := (		
		"00001000000000000000", -- 0		1       	2	_	_	_	
		"00001000010001000011", -- 1		2      	_	_	3	4
		"00011001000010100110", -- 10		3			4	5	6	7
		"00011000110001100010", -- 11		4			_	_	_	3		
		"00101000110001000001", -- 100	5			6	4	3	2		
		"00110000100011000100", -- 101	6			7	3	7	5		
		"11111001010010000011", -- 110	7			32	6	5	4
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000"
	);

BEGIN
	-- saida da memoria
	dado_saida <= memoria(to_integer(unsigned(endereco)));

END ARCHITECTURE rom_modelsim;