LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		enderecoA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		enderecoB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saidaA : OUT STD_LOGIC_VECTOR(27 DOWNTO 0);
		dado_saidaB : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE t_mem IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(27 DOWNTO 0);

	CONSTANT mem : t_mem := (
		-- "1111100000110000100110000110", -- Grafo quebrado
		-- "0000100000000000101010001110",
		-- "0010001001011000000110011010",
		-- "0001100000010000011000000010",
		-- "0000001001000000010110010100",
		-- "0010100000101000001010010000",
		-- "0100101000100000110000011110",
		-- "0101001001100000111000100010",
		-- "0100110001110001001110100100",
		-- "0100001010001100110110100000",
		-- "0110000010111000111110111010",
		-- "0111101010101001011001011100",
		-- "0110101011000001101110101011",
		-- "0110001011010001100110110100",
		-- "1000001010100001110000111000",
		-- "1001101100011001011111000100",
		-- "1001001100101001110111001000",
		-- "1000100011111010001000111100",
		-- "1010001100001010000111000000",
		-- "1010101100110001111111001100",
		-- "1010000101100010010111011010",
		-- "1010100101010010011111010100",
		-- "1011000101000010110001010010",
		-- "1100001110000011001010101100",
		-- "1100111110000010111111011110",
		-- "1100011110010010111011101000",
		-- "1101101110100011010001100100",
		-- "1110110111000011010111110100",
		-- "1111001111101111111011101110",
		-- "1110100110111111101001101100",
		-- "1110010111100011100111111000",
		-- "1111100111110011100011111100",

		"0000001000000000000110000110", -- Quadriculado
		"0000101000000000001110001010",
		"0010101000010000010110001110",
		"0010001000100000011110001110",
		"0100001001010000011110010010",
		"0011001100000000010110010010",
		"0011101001100000101110011010",
		"0100101101010000110111001010",
		"0100001010000000100110100010",
		"0101001010010000111110111010",
		"0101101010100001001110110010",
		"0101101010110001010110110110",
		"0110101010100001100110110010",
		"0110101010110001100110110110",
		"0111001010010001110110111010",
		"0111101011110010000110111110",
		"0111101100010010000110010110",
		"1001101100010010001111000010",
		"1001001001110010010111001010",
		"1010001100110010001111001110",
		"1011001101000010011111010110",
		"1011101101000010101110011110",
		"1100001101100010100111011010",
		"1100101101110010101111011110",
		"1101001110000010110111100010",
		"1110001110010010111111100110",
		"1101101110100011000111110010",
		"1101101110110011010111101110",
		"1110101110100011001111110010",
		"1110101111010011100111111010",
		"1111001111010011110111111110",
		"1111101111100011111111111110",

		"0001001000110000100110000110", -- Grafo
		"0000100000000000101010001110",
		"0010001001011000000110011010",
		"0001100000010000011000000010",
		"0000001001000000010110010100",
		"0010100000101000001010010000",
		"0100101000100000110000011110",
		"0101001001100000111000100010",
		"0100110001110001001110100100",
		"0100001010001100110110100000",
		"0110000010111000111110111010",
		"0111101010101001011001011100",
		"0110101011000001101110101011",
		"0110001011010001100110110100",
		"1000001010100001110000111000",
		"1001101100011001011111000100",
		"1001001100101001110111001000",
		"1000100011111010001000111100",
		"1010001100001010000111000000",
		"1010101100110001111111001100",
		"1010000101100010010111011010",
		"1010100101010010011111010100",
		"1011000101000010110001010010",
		"1100001110000011001010101100",
		"1100111110000010111111011110",
		"1100011110010010111011101000",
		"1101101110100011010001100100",
		"1110110111000011010111110100",
		"1111001111101111111011101110",
		"1110100110111111101001101100",
		"1110010111100011100111111000",
		"1111100111110011100011111100",

		"0000101000000000000001111101", -- Teste
		"0000100000100000000110001010",
		"0001101000010000011110000110",
		"0001001001111000010110010010",
		"0010000000110000101100010000",
		"0011001001000100110110010100",
		"0010101001110000101110011000",
		"1111011000111001000000011010",
		"1111010010000001000000011101",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011111010001111110001111110",
		"1111100111100000000001111100",

		"0000101000000000000001111101",
		"0000100000100000000110001010",
		"0001101000010000011110000110",
		"0001001001111000010110010010",
		"0010000000110000101100010000",
		"0011001001000100110110010100",
		"0010101001110000101110011000",
		"1111011000111001000000011010",
		"1111010010000001000000011101",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011111010001111110001111110",
		"1111100111100000000001111100"
	);

BEGIN
	-- saida da memoria
	dado_saidaA <= mem(to_integer(unsigned(enderecoA)));
	dado_saidaB <= mem(to_integer(unsigned(enderecoB)));

END ARCHITECTURE rom_modelsim;