LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		enderecoA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		enderecoB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saidaA : OUT STD_LOGIC_VECTOR(27 DOWNTO 0);
		dado_saidaB : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE t_mem IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(27 DOWNTO 0);

	CONSTANT mem : t_mem := (
		"0000110000000000000001111110",
		"0000100000101100000000001001",
		"0001110000011100011000000101",
		"0001010001110100010000010001",
		"0010000000111100101010010000",
		"0011010001001000110000010100",
		"0010110001111100101000011000",
		"1111000000110101000110011001",
		"1111001010000001000000011110",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011100010000011110001111101",
		"1111100111101100000111111100",

		"0000110000000000000001111110",
		"0000100000101100000000001001",
		"0001110000011100011000000101",
		"0001010001110100010000010001",
		"0010000000111100101010010000",
		"0011010001001000110000010100",
		"0010110001111100101000011000",
		"1111000000110101000110011001",
		"1111001010000001000000011110",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011100010000011110001111101",
		"1111100111101100000111111100",

		"0000110000000000000001111110",
		"0000100000101100000000001001",
		"0001110000011100011000000101",
		"0001010001110100010000010001",
		"0010000000111100101010010000",
		"0011010001001000110000010100",
		"0010110001111100101000011000",
		"1111000000110101000110011001",
		"1111001010000001000000011110",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011100010000011110001111101",
		"1111100111101100000111111100",

		"0000110000000000000001111110",
		"0000100000101100000000001001",
		"0001110000011100011000000101",
		"0001010001110100010000010001",
		"0010000000111100101010010000",
		"0011010001001000110000010100",
		"0010110001111100101000011000",
		"1111000000110101000110011001",
		"1111001010000001000000011110",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011100010000011110001111101",
		"1111100111101100000111111100"
	);

BEGIN
	-- saida da memoria
	dado_saidaA <= mem(to_integer(unsigned(enderecoA)));
	dado_saidaB <= mem(to_integer(unsigned(enderecoB)));

END ARCHITECTURE rom_modelsim;