library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_128x20 is
   port (       
       endereco     : in  std_logic_vector(6 downto 0);
       dado_saida   : out std_logic_vector(19 downto 0)
    );
end entity rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
architecture rom_modelsim of rom_128x20 is
  type   arranjo_memoria is array(0 to 127) of std_logic_vector(19 downto 0);
  signal memoria : arranjo_memoria := (
                                        "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000",
													 "00000000000000000000"
													 );
  
begin
  -- saida da memoria
  dado_saida <= memoria(to_integer(unsigned(endereco)));

end architecture rom_modelsim;