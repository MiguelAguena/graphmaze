LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		enderecoA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		enderecoB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saidaA : OUT STD_LOGIC_VECTOR(27 DOWNTO 0);
		dado_saidaB : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE t_mem IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(27 DOWNTO 0);

	CONSTANT mem : t_mem := (
		"0000001000000000000110001010", -- Quadriculado
		"0001101000010000001110010010",
		"0001001000000000010110010110",
		"0011001000110000001110001110",
		"0011101000010000100110100010",
		"0100001000100000101110100110",
		"0101001001100000011110101110",
		"0011101001110000100110011110",
		"0110001001000000101110110110",
		"0110101001010001001110100110",
		"0111001010100000110110101010",
		"0111101001100001011111000010",
		"1000001011000001000110110010",
		"1000101010000001001110110110",
		"1001001011100001010110111010",
		"1001101011110001011110111110",
		"1010001010110001100111010110",
		"1000101100010001101111000110",
		"1011001100100001110111011110",
		"1011101100110001111111001110",
		"1100001101000010000111100110",
		"1010101100000010101111010110",
		"1011001101100010010111011010",
		"1101001100100010011111011110",
		"1101101110000010100111110010",
		"1100101101000011001111100110",
		"1101001110100010111111110110",
		"1101101110110011000111111010",
		"1111001110000011100111110010",
		"1110101110100011101111111110",
		"1111001110110011100111111010",
		"1111101111010011111111111110",

		"0000101000000000000001111101", -- Teste
		"0000100000100000000110001010",
		"0001101000010000011110000110",
		"0001001001111000010110010010",
		"0010000000110000101100010000",
		"0011001001000100110110010100",
		"0010101001110000101110011000",
		"1111011000111001000000011010",
		"1111010010000001000000011101",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011111010001111110001111110",
		"1111100111100000000001111100",

		"0000101000000000000001111101",
		"0000100000100000000110001010",
		"0001101000010000011110000110",
		"0001001001111000010110010010",
		"0010000000110000101100010000",
		"0011001001000100110110010100",
		"0010101001110000101110011000",
		"1111011000111001000000011010",
		"1111010010000001000000011101",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011111010001111110001111110",
		"1111100111100000000001111100",

		"0000101000000000000001111101",
		"0000100000100000000110001010",
		"0001101000010000011110000110",
		"0001001001111000010110010010",
		"0010000000110000101100010000",
		"0011001001000100110110010100",
		"0010101001110000101110011000",
		"1111011000111001000000011010",
		"1111010010000001000000011101",
		"0100100010010001001000100100",
		"0101000010100001010000101000",
		"0101100010110001011000101100",
		"0110000011000001100000110000",
		"0110100011010001101000110100",
		"0111000011100001110000111000",
		"0111100011110001111000111100",
		"1000000100000010000001000000",
		"1000100100010010001001000100",
		"1001000100100010010001001000",
		"1001100100110010011001001100",
		"1010000101000010100001010000",
		"1010100101010010101001010100",
		"1011000101100010110001011000",
		"1011100101110010111001011100",
		"1100000110000011000001100000",
		"1100100110010011001001100100",
		"1101000110100011010001101000",
		"1101100110110011011001101100",
		"1110000111000011100001110000",
		"1110100111010011101001110100",
		"0011111010001111110001111110",
		"1111100111100000000001111100");

BEGIN
	-- saida da memoria
	dado_saidaA <= mem(to_integer(unsigned(enderecoA)));
	dado_saidaB <= mem(to_integer(unsigned(enderecoB)));

END ARCHITECTURE rom_modelsim;