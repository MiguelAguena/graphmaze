LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		enderecoA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		enderecoB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saidaA : OUT STD_LOGIC_VECTOR(27 DOWNTO 0);
		dado_saidaB : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE t_mem IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(27 DOWNTO 0);

	CONSTANT mem : t_mem := (

		"0000001000000000000110000110", -- Quadriculado
		"0000101000000000001110001010",
		"0010101000010000010110001110",
		"0010001000100000011110001110",
		"0100001001010000011110010010",
		"0011001100000000010110010010",
		"0011101001100000101110011010",
		"0100101101010000110111001010",
		"0100001010000000100110100010",
		"0101001010010000111110111010",
		"0101101010100001001110110010",
		"0101101010110001010110110110",
		"0110101010100001100110110010",
		"0110101010110001100110110110",
		"0111001010010001110110111010",
		"0111101011110010000110111110",
		"0111101100010010000110010110",
		"1001101100010010001111000010",
		"1001001001110010010111001010",
		"1010001100110010001111001110",
		"1011001101000010011111010110",
		"1011101101000010101110011110",
		"1100001101100010100111011010",
		"1100101101110010101111011110",
		"1101001110000010110111100010",
		"1110001110010010111111100110",
		"1101101110100011000111110010",
		"1101101110110011010111101110",
		"1110101110100011001111110010",
		"1110101111010011100111111010",
		"1111001111010011110111111110",
		"1111101111100011111111111110",

		"0001001000110000100110000110", -- Grafo
		"0000100000000000101010001110",
		"0010001001011000000110011010",
		"0001100000010000011000000010",
		"0000001001000000010110010100",
		"0010100000101000001010010000",
		"0100101000100000110000011110",
		"0101001001100000111000100010",
		"0100110001110001001110100100",
		"0100001010001100110110100000",
		"0110000010111000111110111010",
		"0111101010101001011001011100",
		"0110101011000001101110101011",
		"0110001011010001100110110100",
		"1000001010100001110000111000",
		"1001101100011001011111000100",
		"1001001100101001110111001000",
		"1000100011111010001000111100",
		"1010001100001010000111000000",
		"1010101100110001111111001100",
		"1010000101100010010111011010",
		"1010100101010010011111010100",
		"1011000101000010110001010010",
		"1100001110000011001010101100",
		"1100111110000010111111011110",
		"1100011110010010111011101000",
		"1101101110100011010001100100",
		"1110110111000011010111110100",
		"1111001111101111111011101110",
		"1110100110111111101001101100",
		"1110010111100011100111111000",
		"1111100111110011100011111100",

		"0001011000000000000000000110", -- Salão
		"0001001000000000011110001100",
		"0000011000100000001110001110",
		"0000101000100000100110000100",
		"0001101010000000101110011010",
		"0010001001010001001110010100",
		"0100010001000000110000011110",
		"0110001001100001010110101101",
		"0110101001101101000000010010",
		"0010101010010001001000100100",
		"0011101010111001011110101100",
		"0101001010101000111000101000",
		"0110000011000000111110110000",
		"0111111011110001000110111010",
		"0111000011010001110000111110",
		"0110111011100010000000110110",
		"1001110100010010011010111101",
		"1010001100100010010011000010",
		"1001111100110010001011000110",
		"1001011100001110000011001010",
		"1010101101000010001111011110",
		"1100101101100010100111010100",
		"1101010101100010110001010110",
		"1100000101000010111001101100",
		"1100000110000011011111011111",
		"1101000110010010101111110010",
		"1110001101101111110111100111",
		"1100001110110011101111011100",
		"1110000110010011010111111000",
		"1101101111111011110011110100",
		"1101001111100011101011110000",
		"1111100111011011111001111100",

		"0000101000000001001110000100", -- Corredor
		"0001001000101000000110000000",
		"0001101000011000001110001110",
		"0010001000100000010110010100",
		"0010101010011000011110011000",
		"0011001010010000100110001100",
		"0100101010001000101110010000",
		"1001101010101001000110101100",
		"0011101001101001010110101000",
		"0000001001001000110110010110",
		"0100001001111001011110100000",
		"0101001011001001101110011100",
		"0110000010111001100000111010",
		"0101101100111001111110111100",
		"1000001011000010010001010000",
		"0110101100010010001110110100",
		"1000000100000001110111000000",
		"0111101100110010011110111110",
		"1010101100100010111010111001",
		"1000101011011000111111000110",
		"1010000101110010100000111000",
		"1011001101111010010111011000",
		"1100001101100010101111010100",
		"1011100101011010010011010010",
		"1100101110110010110111110000",
		"1110010110111011000111101010",
		"1110001110010011010001101000",
		"1101100110011011011001100010",
		"1110100110011111010111100000",
		"1111001111010011111111110011",
		"1111000111100011101111111000",
		"1110101111110011111001111100"
	);

BEGIN
	-- saida da memoria
	dado_saidaA <= mem(to_integer(unsigned(enderecoA)));
	dado_saidaB <= mem(to_integer(unsigned(enderecoB)));

END ARCHITECTURE rom_modelsim;