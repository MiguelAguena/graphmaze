LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom_128x20 IS
	PORT (
		enderecoA : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		enderecoB : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dado_saidaA : OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		dado_saidaB : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
	);
END ENTITY rom_128x20;

-- Dados iniciais (para simulacao com Modelsim) 
ARCHITECTURE rom_modelsim OF rom_128x20 IS
	TYPE arranjo_memoria IS ARRAY(0 TO 127) OF STD_LOGIC_VECTOR(19 DOWNTO 0);
	
	-- para ganhar: R L D R
															    --	R	U	L	D
	SIGNAL memoria : arranjo_memoria := (		
		"00001000000000011111", -- 00000			1       	2	_	_	_	
		"00001000010001000011", -- 00001			2      	_	_	3	4
		"00011001000010100110", -- 00010			3			4	5	6	7
		"00011000110001100010", -- 00011			4			_	_	_	3		
		"00101000110001000001", -- 00100		   5			6	4	3	2		
		"00110000100011000100", -- 00101		   6			7	3	7	5		
		"11110001010010000011", -- 00110		   7			31	6	5	4
		"00000000000000000000", -- 00111
		"00000000000000000000", -- 01000
		"00000000000000000000", -- 01001
		"00000000000000000000", -- 01010
		"00000000000000000000", -- 01011
		"00000000000000000000", -- 01100
		"00000000000000000000", -- 01101
		"00000000000000000000", -- 01110
		"00000000000000000000", -- 01111
		"00000000000000000000", -- 10000
		"00000000000000000000", -- 10001
		"00000000000000000000", -- 10010
		"00000000000000000000", -- 10011
		"00000000000000000000", -- 10100
		"00000000000000000000", -- 10101
		"00000000000000000000", -- 10110
		"00000000000000000000", -- 10111
		"00000000000000000000", -- 11000
		"00000000000000000000", -- 11001
		"00000000000000000000", -- 11010
		"00000000000000000000", -- 11011
		"00000000000000000000", -- 11100
		"00000000000000000000", -- 11101
		"00110001100011011111", -- 11110		   31			7	7	7	32
		"11110111101111011110", -- 11111
		"00001000000000000000",
		"00010000000000000000",
		"00011000000000000000",
		"00100000000000000000",
		"00101000000000000000",
		"00110000000000000000",
		"00111000000000000000",
		"01000000000000000000",
		"01001000000000000000",
		"01010000000000000000",
		"01011000000000000000",
		"01100000000000000000",
		"01101000000000000000",
		"01110000000000000000",
		"01111000000000000000",
		"10000000000000000000",
		"10001000000000000000",
		"10010000000000000000",
		"10011000000000000000",
		"10100000000000000000",
		"10101000000000000000",
		"10110000000000000000",
		"10111000000000000000",
		"11000000000000000000",
		"11001000000000000000",
		"11010000000000000000",
		"11011000000000000000",
		"11100000000000000000",
		"11101000000000000000",
		"11110000000000000000",
		"11111000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000",
		"00000000000000000000"
	);

BEGIN
	-- saida da memoria
	dado_saidaA <= memoria(to_integer(unsigned(enderecoA)));
	dado_saidaB <= memoria(to_integer(unsigned(enderecoB)));

END ARCHITECTURE rom_modelsim;